`ifndef BLOCK_EA_VH
`define BLOCK_EA_VH
`define BLOCK_EA_VERSION_BIT_WIDTH 32
`define BLOCK_EA_VERSION_BIT_MASK 32'hffffffff
`define BLOCK_EA_VERSION_BIT_OFFSET 0
`define BLOCK_EA_VERSION_BYTE_WIDTH 4
`define BLOCK_EA_VERSION_BYTE_SIZE 4
`define BLOCK_EA_VERSION_BYTE_OFFSET 10'h000
`define BLOCK_EA_RESET_BIT_WIDTH 32
`define BLOCK_EA_RESET_BIT_MASK 32'hffffffff
`define BLOCK_EA_RESET_BIT_OFFSET 0
`define BLOCK_EA_RESET_BYTE_WIDTH 4
`define BLOCK_EA_RESET_BYTE_SIZE 4
`define BLOCK_EA_RESET_BYTE_OFFSET 10'h00c
`define BLOCK_EA_INDEX_BIT_WIDTH 32
`define BLOCK_EA_INDEX_BIT_MASK 32'hffffffff
`define BLOCK_EA_INDEX_BIT_OFFSET 0
`define BLOCK_EA_INDEX_BYTE_WIDTH 4
`define BLOCK_EA_INDEX_BYTE_SIZE 4
`define BLOCK_EA_INDEX_BYTE_OFFSET 10'h010
`define BLOCK_EA_UART_BIT_RATE_BIT_WIDTH 32
`define BLOCK_EA_UART_BIT_RATE_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_BIT_RATE_BIT_OFFSET 0
`define BLOCK_EA_UART_BIT_RATE_BYTE_WIDTH 4
`define BLOCK_EA_UART_BIT_RATE_BYTE_SIZE 4
`define BLOCK_EA_UART_BIT_RATE_BYTE_OFFSET 10'h100
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BYTE_OFFSET 10'h104
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BYTE_OFFSET 10'h108
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BYTE_OFFSET 10'h10c
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BYTE_OFFSET 10'h110
`define BLOCK_EA_UART_RECV_DATA_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_RECV_DATA_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_RECV_DATA_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_RECV_DATA_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_RECV_DATA_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_RECV_DATA_COUNT_BYTE_OFFSET 10'h114
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BIT_WIDTH 32
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BIT_OFFSET 0
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BYTE_WIDTH 4
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BYTE_SIZE 4
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BYTE_OFFSET 10'h120
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BIT_WIDTH 32
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BIT_OFFSET 0
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BYTE_WIDTH 4
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BYTE_SIZE 4
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BYTE_OFFSET 10'h124
`define BLOCK_EA_MAC_SEND_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_SEND_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_SEND_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_SEND_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_SEND_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_SEND_COUNT_BYTE_OFFSET 10'h200
`define BLOCK_EA_MAC_RECV_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_RECV_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_RECV_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_RECV_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_RECV_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_RECV_COUNT_BYTE_OFFSET 10'h204
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BYTE_OFFSET 10'h210
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BYTE_OFFSET 10'h214
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BYTE_OFFSET 10'h218
`endif
