`ifndef __HEAD_VH__
`define __HEAD_VH__

`define DO_DPA
`define IS_CLIENT
`define VERSION 32'h24072300
`define UART_BITS 8

`endif // __HEAD_VH__