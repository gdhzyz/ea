`ifndef __HEAD_VH__
`define __HEAD_VH__

//`define DO_DPA
//`define DO_DPA_INSIDE_MAC
`define IS_CLIENT
`define VERSION 32'h24072300
`define UART_BITS 8
`define I2S_IN

`endif // __HEAD_VH__