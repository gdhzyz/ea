
`define IS_CLIENT