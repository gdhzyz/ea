package block_ea_rtl_pkg;
  localparam int VERSION_BYTE_WIDTH = 4;
  localparam int VERSION_BYTE_SIZE = 4;
  localparam bit [15:0] VERSION_BYTE_OFFSET = 16'h0000;
  localparam int VERSION_BIT_WIDTH = 32;
  localparam bit [31:0] VERSION_BIT_MASK = 32'hffffffff;
  localparam int VERSION_BIT_OFFSET = 0;
  localparam int RESET_BYTE_WIDTH = 4;
  localparam int RESET_BYTE_SIZE = 4;
  localparam bit [15:0] RESET_BYTE_OFFSET = 16'h000c;
  localparam int RESET_BIT_WIDTH = 1;
  localparam bit RESET_BIT_MASK = 1'h1;
  localparam int RESET_BIT_OFFSET = 0;
  localparam int INDEX_BYTE_WIDTH = 4;
  localparam int INDEX_BYTE_SIZE = 4;
  localparam bit [15:0] INDEX_BYTE_OFFSET = 16'h0010;
  localparam int INDEX_BIT_WIDTH = 4;
  localparam bit [3:0] INDEX_BIT_MASK = 4'hf;
  localparam int INDEX_BIT_OFFSET = 0;
  localparam int UART_BIT_RATE_BYTE_WIDTH = 4;
  localparam int UART_BIT_RATE_BYTE_SIZE = 4;
  localparam bit [15:0] UART_BIT_RATE_BYTE_OFFSET = 16'h0100;
  localparam int UART_BIT_RATE_BIT_WIDTH = 17;
  localparam bit [16:0] UART_BIT_RATE_BIT_MASK = 17'h1ffff;
  localparam int UART_BIT_RATE_BIT_OFFSET = 0;
  localparam int UART_REG_WRITE_REQ_COUNT_BYTE_WIDTH = 4;
  localparam int UART_REG_WRITE_REQ_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] UART_REG_WRITE_REQ_COUNT_BYTE_OFFSET = 16'h0104;
  localparam int UART_REG_WRITE_REQ_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] UART_REG_WRITE_REQ_COUNT_BIT_MASK = 32'hffffffff;
  localparam int UART_REG_WRITE_REQ_COUNT_BIT_OFFSET = 0;
  localparam int UART_REG_READ_REQ_COUNT_BYTE_WIDTH = 4;
  localparam int UART_REG_READ_REQ_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] UART_REG_READ_REQ_COUNT_BYTE_OFFSET = 16'h0108;
  localparam int UART_REG_READ_REQ_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] UART_REG_READ_REQ_COUNT_BIT_MASK = 32'hffffffff;
  localparam int UART_REG_READ_REQ_COUNT_BIT_OFFSET = 0;
  localparam int UART_REG_READ_ACK_COUNT_BYTE_WIDTH = 4;
  localparam int UART_REG_READ_ACK_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] UART_REG_READ_ACK_COUNT_BYTE_OFFSET = 16'h010c;
  localparam int UART_REG_READ_ACK_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] UART_REG_READ_ACK_COUNT_BIT_MASK = 32'hffffffff;
  localparam int UART_REG_READ_ACK_COUNT_BIT_OFFSET = 0;
  localparam int UART_WRITE_DATA_COUNT_BYTE_WIDTH = 4;
  localparam int UART_WRITE_DATA_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] UART_WRITE_DATA_COUNT_BYTE_OFFSET = 16'h0110;
  localparam int UART_WRITE_DATA_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] UART_WRITE_DATA_COUNT_BIT_MASK = 32'hffffffff;
  localparam int UART_WRITE_DATA_COUNT_BIT_OFFSET = 0;
  localparam int UART_RECV_DATA_COUNT_BYTE_WIDTH = 4;
  localparam int UART_RECV_DATA_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] UART_RECV_DATA_COUNT_BYTE_OFFSET = 16'h0114;
  localparam int UART_RECV_DATA_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] UART_RECV_DATA_COUNT_BIT_MASK = 32'hffffffff;
  localparam int UART_RECV_DATA_COUNT_BIT_OFFSET = 0;
  localparam int UART_DATA_DST_FPGA_INDEX_BYTE_WIDTH = 4;
  localparam int UART_DATA_DST_FPGA_INDEX_BYTE_SIZE = 4;
  localparam bit [15:0] UART_DATA_DST_FPGA_INDEX_BYTE_OFFSET = 16'h0120;
  localparam int UART_DATA_DST_FPGA_INDEX_BIT_WIDTH = 4;
  localparam bit [3:0] UART_DATA_DST_FPGA_INDEX_BIT_MASK = 4'hf;
  localparam int UART_DATA_DST_FPGA_INDEX_BIT_OFFSET = 0;
  localparam int UART_REG_DST_FPGA_INDEX_BYTE_WIDTH = 4;
  localparam int UART_REG_DST_FPGA_INDEX_BYTE_SIZE = 4;
  localparam bit [15:0] UART_REG_DST_FPGA_INDEX_BYTE_OFFSET = 16'h0124;
  localparam int UART_REG_DST_FPGA_INDEX_BIT_WIDTH = 4;
  localparam bit [3:0] UART_REG_DST_FPGA_INDEX_BIT_MASK = 4'hf;
  localparam int UART_REG_DST_FPGA_INDEX_BIT_OFFSET = 0;
  localparam int MAC_SEND_COUNT_BYTE_WIDTH = 4;
  localparam int MAC_SEND_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_SEND_COUNT_BYTE_OFFSET = 16'h0200;
  localparam int MAC_SEND_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] MAC_SEND_COUNT_BIT_MASK = 32'hffffffff;
  localparam int MAC_SEND_COUNT_BIT_OFFSET = 0;
  localparam int MAC_RECV_COUNT_BYTE_WIDTH = 4;
  localparam int MAC_RECV_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_RECV_COUNT_BYTE_OFFSET = 16'h0204;
  localparam int MAC_RECV_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] MAC_RECV_COUNT_BIT_MASK = 32'hffffffff;
  localparam int MAC_RECV_COUNT_BIT_OFFSET = 0;
  localparam int MAC_REG_WRITE_REQ_COUNT_BYTE_WIDTH = 4;
  localparam int MAC_REG_WRITE_REQ_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_REG_WRITE_REQ_COUNT_BYTE_OFFSET = 16'h0210;
  localparam int MAC_REG_WRITE_REQ_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] MAC_REG_WRITE_REQ_COUNT_BIT_MASK = 32'hffffffff;
  localparam int MAC_REG_WRITE_REQ_COUNT_BIT_OFFSET = 0;
  localparam int MAC_REG_READ_REQ_COUNT_BYTE_WIDTH = 4;
  localparam int MAC_REG_READ_REQ_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_REG_READ_REQ_COUNT_BYTE_OFFSET = 16'h0214;
  localparam int MAC_REG_READ_REQ_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] MAC_REG_READ_REQ_COUNT_BIT_MASK = 32'hffffffff;
  localparam int MAC_REG_READ_REQ_COUNT_BIT_OFFSET = 0;
  localparam int MAC_REG_READ_ACK_COUNT_BYTE_WIDTH = 4;
  localparam int MAC_REG_READ_ACK_COUNT_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_REG_READ_ACK_COUNT_BYTE_OFFSET = 16'h0218;
  localparam int MAC_REG_READ_ACK_COUNT_BIT_WIDTH = 32;
  localparam bit [31:0] MAC_REG_READ_ACK_COUNT_BIT_MASK = 32'hffffffff;
  localparam int MAC_REG_READ_ACK_COUNT_BIT_OFFSET = 0;
  localparam int MAC_DLY_SEL_BYTE_WIDTH = 4;
  localparam int MAC_DLY_SEL_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_DLY_SEL_BYTE_OFFSET = 16'h0300;
  localparam int MAC_DLY_SEL_BIT_WIDTH = 3;
  localparam bit [2:0] MAC_DLY_SEL_BIT_MASK = 3'h7;
  localparam int MAC_DLY_SEL_BIT_OFFSET = 0;
  localparam int MAC_DLY_INC_BYTE_WIDTH = 4;
  localparam int MAC_DLY_INC_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_DLY_INC_BYTE_OFFSET = 16'h0304;
  localparam int MAC_DLY_INC_BIT_WIDTH = 1;
  localparam bit MAC_DLY_INC_BIT_MASK = 1'h1;
  localparam int MAC_DLY_INC_BIT_OFFSET = 0;
  localparam int MAC_DLY_VALUE_BYTE_WIDTH = 4;
  localparam int MAC_DLY_VALUE_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_DLY_VALUE_BYTE_OFFSET = 16'h0308;
  localparam int MAC_DLY_VALUE_BIT_WIDTH = 5;
  localparam bit [4:0] MAC_DLY_VALUE_BIT_MASK = 5'h1f;
  localparam int MAC_DLY_VALUE_BIT_OFFSET = 0;
  localparam int MAC_ENABLE_JUMBO_TEST_BYTE_WIDTH = 4;
  localparam int MAC_ENABLE_JUMBO_TEST_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_ENABLE_JUMBO_TEST_BYTE_OFFSET = 16'h030c;
  localparam int MAC_ENABLE_JUMBO_TEST_BIT_WIDTH = 1;
  localparam bit MAC_ENABLE_JUMBO_TEST_BIT_MASK = 1'h1;
  localparam int MAC_ENABLE_JUMBO_TEST_BIT_OFFSET = 0;
  localparam int MAC_JUMBO_ERROR_BYTE_WIDTH = 4;
  localparam int MAC_JUMBO_ERROR_BYTE_SIZE = 4;
  localparam bit [15:0] MAC_JUMBO_ERROR_BYTE_OFFSET = 16'h0310;
  localparam int MAC_JUMBO_ERROR_BIT_WIDTH = 1;
  localparam bit MAC_JUMBO_ERROR_BIT_MASK = 1'h1;
  localparam int MAC_JUMBO_ERROR_BIT_OFFSET = 0;
  localparam int MAC_TEST_ARRAY_BYTE_WIDTH = 64;
  localparam int MAC_TEST_ARRAY_BYTE_SIZE = 64;
  localparam bit [15:0] MAC_TEST_ARRAY_BYTE_OFFSET = 16'h0400;
  localparam int MAC_TEST_ARRAY_BIT_WIDTH = 32;
  localparam bit [31:0] MAC_TEST_ARRAY_BIT_MASK = 32'hffffffff;
  localparam int MAC_TEST_ARRAY_BIT_OFFSET[16] = '{0, 32, 64, 96, 128, 160, 192, 224, 256, 288, 320, 352, 384, 416, 448, 480};
  localparam int I2S_OUT_TDM_NUM_BYTE_WIDTH = 16;
  localparam int I2S_OUT_TDM_NUM_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_TDM_NUM_BYTE_OFFSET = 16'h1000;
  localparam int I2S_OUT_TDM_NUM_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_TDM_NUM_BIT_MASK = 8'hff;
  localparam int I2S_OUT_TDM_NUM_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_IS_MASTER_BYTE_WIDTH = 16;
  localparam int I2S_OUT_IS_MASTER_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_IS_MASTER_BYTE_OFFSET = 16'h1010;
  localparam int I2S_OUT_IS_MASTER_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_IS_MASTER_BIT_MASK = 8'hff;
  localparam int I2S_OUT_IS_MASTER_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_ENABLE_BYTE_WIDTH = 16;
  localparam int I2S_OUT_ENABLE_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_ENABLE_BYTE_OFFSET = 16'h1020;
  localparam int I2S_OUT_ENABLE_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_ENABLE_BIT_MASK = 8'hff;
  localparam int I2S_OUT_ENABLE_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_FPGA_INDEX_BYTE_WIDTH = 16;
  localparam int I2S_OUT_FPGA_INDEX_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_FPGA_INDEX_BYTE_OFFSET = 16'h1030;
  localparam int I2S_OUT_FPGA_INDEX_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_FPGA_INDEX_BIT_MASK = 8'hff;
  localparam int I2S_OUT_FPGA_INDEX_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_WORD_WIDTH_BYTE_WIDTH = 16;
  localparam int I2S_OUT_WORD_WIDTH_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_WORD_WIDTH_BYTE_OFFSET = 16'h1040;
  localparam int I2S_OUT_WORD_WIDTH_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_WORD_WIDTH_BIT_MASK = 8'hff;
  localparam int I2S_OUT_WORD_WIDTH_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_VALID_WORD_WIDTH_BYTE_WIDTH = 16;
  localparam int I2S_OUT_VALID_WORD_WIDTH_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_VALID_WORD_WIDTH_BYTE_OFFSET = 16'h1050;
  localparam int I2S_OUT_VALID_WORD_WIDTH_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_VALID_WORD_WIDTH_BIT_MASK = 8'hff;
  localparam int I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_LRCK_IS_PULSE_BYTE_WIDTH = 16;
  localparam int I2S_OUT_LRCK_IS_PULSE_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_LRCK_IS_PULSE_BYTE_OFFSET = 16'h1060;
  localparam int I2S_OUT_LRCK_IS_PULSE_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_LRCK_IS_PULSE_BIT_MASK = 8'hff;
  localparam int I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_LRCK_POLARITY_BYTE_WIDTH = 16;
  localparam int I2S_OUT_LRCK_POLARITY_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_LRCK_POLARITY_BYTE_OFFSET = 16'h1070;
  localparam int I2S_OUT_LRCK_POLARITY_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_LRCK_POLARITY_BIT_MASK = 8'hff;
  localparam int I2S_OUT_LRCK_POLARITY_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_LRCK_ALIGNMENT_BYTE_WIDTH = 16;
  localparam int I2S_OUT_LRCK_ALIGNMENT_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_LRCK_ALIGNMENT_BYTE_OFFSET = 16'h1080;
  localparam int I2S_OUT_LRCK_ALIGNMENT_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_LRCK_ALIGNMENT_BIT_MASK = 8'hff;
  localparam int I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_I2S_INDEX_BYTE_WIDTH = 16;
  localparam int I2S_OUT_I2S_INDEX_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_OUT_I2S_INDEX_BYTE_OFFSET = 16'h1090;
  localparam int I2S_OUT_I2S_INDEX_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_OUT_I2S_INDEX_BIT_MASK = 8'hff;
  localparam int I2S_OUT_I2S_INDEX_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_OUT_FRAME_NUM_BYTE_WIDTH = 64;
  localparam int I2S_OUT_FRAME_NUM_BYTE_SIZE = 64;
  localparam bit [15:0] I2S_OUT_FRAME_NUM_BYTE_OFFSET = 16'h1100;
  localparam int I2S_OUT_FRAME_NUM_BIT_WIDTH = 32;
  localparam bit [31:0] I2S_OUT_FRAME_NUM_BIT_MASK = 32'hffffffff;
  localparam int I2S_OUT_FRAME_NUM_BIT_OFFSET[16] = '{0, 32, 64, 96, 128, 160, 192, 224, 256, 288, 320, 352, 384, 416, 448, 480};
  localparam int I2S_OUT_BCLK_FREQ_BYTE_WIDTH = 64;
  localparam int I2S_OUT_BCLK_FREQ_BYTE_SIZE = 64;
  localparam bit [15:0] I2S_OUT_BCLK_FREQ_BYTE_OFFSET = 16'h1300;
  localparam int I2S_OUT_BCLK_FREQ_BIT_WIDTH = 32;
  localparam bit [31:0] I2S_OUT_BCLK_FREQ_BIT_MASK = 32'hffffffff;
  localparam int I2S_OUT_BCLK_FREQ_BIT_OFFSET[16] = '{0, 32, 64, 96, 128, 160, 192, 224, 256, 288, 320, 352, 384, 416, 448, 480};
  localparam int I2S_IN_TDM_NUM_BYTE_WIDTH = 16;
  localparam int I2S_IN_TDM_NUM_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_TDM_NUM_BYTE_OFFSET = 16'h4000;
  localparam int I2S_IN_TDM_NUM_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_TDM_NUM_BIT_MASK = 8'hff;
  localparam int I2S_IN_TDM_NUM_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_IS_MASTER_BYTE_WIDTH = 16;
  localparam int I2S_IN_IS_MASTER_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_IS_MASTER_BYTE_OFFSET = 16'h4010;
  localparam int I2S_IN_IS_MASTER_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_IS_MASTER_BIT_MASK = 8'hff;
  localparam int I2S_IN_IS_MASTER_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_ENABLE_BYTE_WIDTH = 16;
  localparam int I2S_IN_ENABLE_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_ENABLE_BYTE_OFFSET = 16'h4020;
  localparam int I2S_IN_ENABLE_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_ENABLE_BIT_MASK = 8'hff;
  localparam int I2S_IN_ENABLE_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_FPGA_INDEX_BYTE_WIDTH = 16;
  localparam int I2S_IN_FPGA_INDEX_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_FPGA_INDEX_BYTE_OFFSET = 16'h4030;
  localparam int I2S_IN_FPGA_INDEX_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_FPGA_INDEX_BIT_MASK = 8'hff;
  localparam int I2S_IN_FPGA_INDEX_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_WORD_WIDTH_BYTE_WIDTH = 16;
  localparam int I2S_IN_WORD_WIDTH_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_WORD_WIDTH_BYTE_OFFSET = 16'h4040;
  localparam int I2S_IN_WORD_WIDTH_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_WORD_WIDTH_BIT_MASK = 8'hff;
  localparam int I2S_IN_WORD_WIDTH_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_VALID_WORD_WIDTH_BYTE_WIDTH = 16;
  localparam int I2S_IN_VALID_WORD_WIDTH_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_VALID_WORD_WIDTH_BYTE_OFFSET = 16'h4050;
  localparam int I2S_IN_VALID_WORD_WIDTH_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_VALID_WORD_WIDTH_BIT_MASK = 8'hff;
  localparam int I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_LRCK_IS_PULSE_BYTE_WIDTH = 16;
  localparam int I2S_IN_LRCK_IS_PULSE_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_LRCK_IS_PULSE_BYTE_OFFSET = 16'h4060;
  localparam int I2S_IN_LRCK_IS_PULSE_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_LRCK_IS_PULSE_BIT_MASK = 8'hff;
  localparam int I2S_IN_LRCK_IS_PULSE_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_LRCK_POLARITY_BYTE_WIDTH = 16;
  localparam int I2S_IN_LRCK_POLARITY_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_LRCK_POLARITY_BYTE_OFFSET = 16'h4070;
  localparam int I2S_IN_LRCK_POLARITY_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_LRCK_POLARITY_BIT_MASK = 8'hff;
  localparam int I2S_IN_LRCK_POLARITY_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_LRCK_ALIGNMENT_BYTE_WIDTH = 16;
  localparam int I2S_IN_LRCK_ALIGNMENT_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_LRCK_ALIGNMENT_BYTE_OFFSET = 16'h4080;
  localparam int I2S_IN_LRCK_ALIGNMENT_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_LRCK_ALIGNMENT_BIT_MASK = 8'hff;
  localparam int I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_I2S_INDEX_BYTE_WIDTH = 16;
  localparam int I2S_IN_I2S_INDEX_BYTE_SIZE = 16;
  localparam bit [15:0] I2S_IN_I2S_INDEX_BYTE_OFFSET = 16'h4090;
  localparam int I2S_IN_I2S_INDEX_BIT_WIDTH = 8;
  localparam bit [7:0] I2S_IN_I2S_INDEX_BIT_MASK = 8'hff;
  localparam int I2S_IN_I2S_INDEX_BIT_OFFSET[16] = '{0, 8, 16, 24, 32, 40, 48, 56, 64, 72, 80, 88, 96, 104, 112, 120};
  localparam int I2S_IN_FRAME_NUM_BYTE_WIDTH = 64;
  localparam int I2S_IN_FRAME_NUM_BYTE_SIZE = 64;
  localparam bit [15:0] I2S_IN_FRAME_NUM_BYTE_OFFSET = 16'h4100;
  localparam int I2S_IN_FRAME_NUM_BIT_WIDTH = 32;
  localparam bit [31:0] I2S_IN_FRAME_NUM_BIT_MASK = 32'hffffffff;
  localparam int I2S_IN_FRAME_NUM_BIT_OFFSET[16] = '{0, 32, 64, 96, 128, 160, 192, 224, 256, 288, 320, 352, 384, 416, 448, 480};
  localparam int I2S_IN_BCLK_FREQ_BYTE_WIDTH = 64;
  localparam int I2S_IN_BCLK_FREQ_BYTE_SIZE = 64;
  localparam bit [15:0] I2S_IN_BCLK_FREQ_BYTE_OFFSET = 16'h4300;
  localparam int I2S_IN_BCLK_FREQ_BIT_WIDTH = 32;
  localparam bit [31:0] I2S_IN_BCLK_FREQ_BIT_MASK = 32'hffffffff;
  localparam int I2S_IN_BCLK_FREQ_BIT_OFFSET[16] = '{0, 32, 64, 96, 128, 160, 192, 224, 256, 288, 320, 352, 384, 416, 448, 480};
endpackage
