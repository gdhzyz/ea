`ifndef BLOCK_EA_VH
`define BLOCK_EA_VH
`define BLOCK_EA_VERSION_BIT_WIDTH 32
`define BLOCK_EA_VERSION_BIT_MASK 32'hffffffff
`define BLOCK_EA_VERSION_BIT_OFFSET 0
`define BLOCK_EA_VERSION_BYTE_WIDTH 4
`define BLOCK_EA_VERSION_BYTE_SIZE 4
`define BLOCK_EA_VERSION_BYTE_OFFSET 16'h0000
`define BLOCK_EA_RESET_BIT_WIDTH 1
`define BLOCK_EA_RESET_BIT_MASK 1'h1
`define BLOCK_EA_RESET_BIT_OFFSET 0
`define BLOCK_EA_RESET_BYTE_WIDTH 4
`define BLOCK_EA_RESET_BYTE_SIZE 4
`define BLOCK_EA_RESET_BYTE_OFFSET 16'h000c
`define BLOCK_EA_INDEX_BIT_WIDTH 4
`define BLOCK_EA_INDEX_BIT_MASK 4'hf
`define BLOCK_EA_INDEX_BIT_OFFSET 0
`define BLOCK_EA_INDEX_BYTE_WIDTH 4
`define BLOCK_EA_INDEX_BYTE_SIZE 4
`define BLOCK_EA_INDEX_BYTE_OFFSET 16'h0010
`define BLOCK_EA_UART_BIT_RATE_BIT_WIDTH 17
`define BLOCK_EA_UART_BIT_RATE_BIT_MASK 17'h1ffff
`define BLOCK_EA_UART_BIT_RATE_BIT_OFFSET 0
`define BLOCK_EA_UART_BIT_RATE_BYTE_WIDTH 4
`define BLOCK_EA_UART_BIT_RATE_BYTE_SIZE 4
`define BLOCK_EA_UART_BIT_RATE_BYTE_OFFSET 16'h0100
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_REG_WRITE_REQ_COUNT_BYTE_OFFSET 16'h0104
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_REG_READ_REQ_COUNT_BYTE_OFFSET 16'h0108
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_REG_READ_ACK_COUNT_BYTE_OFFSET 16'h010c
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_WRITE_DATA_COUNT_BYTE_OFFSET 16'h0110
`define BLOCK_EA_UART_RECV_DATA_COUNT_BIT_WIDTH 32
`define BLOCK_EA_UART_RECV_DATA_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_UART_RECV_DATA_COUNT_BIT_OFFSET 0
`define BLOCK_EA_UART_RECV_DATA_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_UART_RECV_DATA_COUNT_BYTE_SIZE 4
`define BLOCK_EA_UART_RECV_DATA_COUNT_BYTE_OFFSET 16'h0114
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BIT_WIDTH 4
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BIT_MASK 4'hf
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BIT_OFFSET 0
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BYTE_WIDTH 4
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BYTE_SIZE 4
`define BLOCK_EA_UART_DATA_DST_FPGA_INDEX_BYTE_OFFSET 16'h0120
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BIT_WIDTH 4
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BIT_MASK 4'hf
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BIT_OFFSET 0
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BYTE_WIDTH 4
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BYTE_SIZE 4
`define BLOCK_EA_UART_REG_DST_FPGA_INDEX_BYTE_OFFSET 16'h0124
`define BLOCK_EA_MAC_SEND_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_SEND_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_SEND_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_SEND_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_SEND_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_SEND_COUNT_BYTE_OFFSET 16'h0200
`define BLOCK_EA_MAC_RECV_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_RECV_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_RECV_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_RECV_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_RECV_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_RECV_COUNT_BYTE_OFFSET 16'h0204
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_REG_WRITE_REQ_COUNT_BYTE_OFFSET 16'h0210
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_REG_READ_REQ_COUNT_BYTE_OFFSET 16'h0214
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BIT_WIDTH 32
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BIT_OFFSET 0
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BYTE_WIDTH 4
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BYTE_SIZE 4
`define BLOCK_EA_MAC_REG_READ_ACK_COUNT_BYTE_OFFSET 16'h0218
`define BLOCK_EA_MAC_DLY_SEL_BIT_WIDTH 3
`define BLOCK_EA_MAC_DLY_SEL_BIT_MASK 3'h7
`define BLOCK_EA_MAC_DLY_SEL_BIT_OFFSET 0
`define BLOCK_EA_MAC_DLY_SEL_BYTE_WIDTH 4
`define BLOCK_EA_MAC_DLY_SEL_BYTE_SIZE 4
`define BLOCK_EA_MAC_DLY_SEL_BYTE_OFFSET 16'h0300
`define BLOCK_EA_MAC_DLY_INC_BIT_WIDTH 1
`define BLOCK_EA_MAC_DLY_INC_BIT_MASK 1'h1
`define BLOCK_EA_MAC_DLY_INC_BIT_OFFSET 0
`define BLOCK_EA_MAC_DLY_INC_BYTE_WIDTH 4
`define BLOCK_EA_MAC_DLY_INC_BYTE_SIZE 4
`define BLOCK_EA_MAC_DLY_INC_BYTE_OFFSET 16'h0304
`define BLOCK_EA_MAC_DLY_VALUE_BIT_WIDTH 5
`define BLOCK_EA_MAC_DLY_VALUE_BIT_MASK 5'h1f
`define BLOCK_EA_MAC_DLY_VALUE_BIT_OFFSET 0
`define BLOCK_EA_MAC_DLY_VALUE_BYTE_WIDTH 4
`define BLOCK_EA_MAC_DLY_VALUE_BYTE_SIZE 4
`define BLOCK_EA_MAC_DLY_VALUE_BYTE_OFFSET 16'h0308
`define BLOCK_EA_MAC_ENABLE_JUMBO_TEST_BIT_WIDTH 1
`define BLOCK_EA_MAC_ENABLE_JUMBO_TEST_BIT_MASK 1'h1
`define BLOCK_EA_MAC_ENABLE_JUMBO_TEST_BIT_OFFSET 0
`define BLOCK_EA_MAC_ENABLE_JUMBO_TEST_BYTE_WIDTH 4
`define BLOCK_EA_MAC_ENABLE_JUMBO_TEST_BYTE_SIZE 4
`define BLOCK_EA_MAC_ENABLE_JUMBO_TEST_BYTE_OFFSET 16'h030c
`define BLOCK_EA_MAC_JUMBO_ERROR_BIT_WIDTH 1
`define BLOCK_EA_MAC_JUMBO_ERROR_BIT_MASK 1'h1
`define BLOCK_EA_MAC_JUMBO_ERROR_BIT_OFFSET 0
`define BLOCK_EA_MAC_JUMBO_ERROR_BYTE_WIDTH 4
`define BLOCK_EA_MAC_JUMBO_ERROR_BYTE_SIZE 4
`define BLOCK_EA_MAC_JUMBO_ERROR_BYTE_OFFSET 16'h0310
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_WIDTH 32
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_MASK 32'hffffffff
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_0 0
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_1 32
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_2 64
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_3 96
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_4 128
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_5 160
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_6 192
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_7 224
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_8 256
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_9 288
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_10 320
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_11 352
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_12 384
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_13 416
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_14 448
`define BLOCK_EA_MAC_TEST_ARRAY_BIT_OFFSET_15 480
`define BLOCK_EA_MAC_TEST_ARRAY_BYTE_WIDTH 64
`define BLOCK_EA_MAC_TEST_ARRAY_BYTE_SIZE 64
`define BLOCK_EA_MAC_TEST_ARRAY_BYTE_OFFSET 16'h0400
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_TDM_NUM_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_TDM_NUM_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_TDM_NUM_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_TDM_NUM_BYTE_OFFSET 16'h1000
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_IS_MASTER_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_IS_MASTER_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_IS_MASTER_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_IS_MASTER_BYTE_OFFSET 16'h1010
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_ENABLE_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_ENABLE_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_ENABLE_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_ENABLE_BYTE_OFFSET 16'h1020
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_FPGA_INDEX_BYTE_OFFSET 16'h1030
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_WORD_WIDTH_BYTE_OFFSET 16'h1040
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_VALID_WORD_WIDTH_BYTE_OFFSET 16'h1050
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_LRCK_IS_PULSE_BYTE_OFFSET 16'h1060
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_LRCK_POLARITY_BYTE_OFFSET 16'h1070
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_LRCK_ALIGNMENT_BYTE_OFFSET 16'h1080
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_WIDTH 8
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_MASK 8'hff
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BYTE_WIDTH 16
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BYTE_SIZE 16
`define BLOCK_EA_I2S_OUT_I2S_INDEX_BYTE_OFFSET 16'h1090
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_WIDTH 32
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_MASK 32'hffffffff
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_1 32
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_2 64
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_3 96
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_4 128
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_5 160
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_6 192
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_7 224
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_8 256
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_9 288
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_10 320
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_11 352
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_12 384
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_13 416
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_14 448
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BIT_OFFSET_15 480
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BYTE_WIDTH 64
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BYTE_SIZE 64
`define BLOCK_EA_I2S_OUT_FRAME_NUM_BYTE_OFFSET 16'h1100
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_WIDTH 32
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_MASK 32'hffffffff
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_1 32
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_2 64
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_3 96
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_4 128
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_5 160
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_6 192
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_7 224
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_8 256
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_9 288
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_10 320
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_11 352
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_12 384
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_13 416
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_14 448
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BIT_OFFSET_15 480
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BYTE_WIDTH 64
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BYTE_SIZE 64
`define BLOCK_EA_I2S_OUT_BCLK_FREQ_BYTE_OFFSET 16'h1300
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_TDM_NUM_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_TDM_NUM_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_TDM_NUM_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_TDM_NUM_BYTE_OFFSET 16'h4000
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_IS_MASTER_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_IS_MASTER_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_IS_MASTER_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_IS_MASTER_BYTE_OFFSET 16'h4010
`define BLOCK_EA_I2S_IN_ENABLE_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_ENABLE_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_ENABLE_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_ENABLE_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_ENABLE_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_ENABLE_BYTE_OFFSET 16'h4020
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_FPGA_INDEX_BYTE_OFFSET 16'h4030
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_WORD_WIDTH_BYTE_OFFSET 16'h4040
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_VALID_WORD_WIDTH_BYTE_OFFSET 16'h4050
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_LRCK_IS_PULSE_BYTE_OFFSET 16'h4060
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_LRCK_POLARITY_BYTE_OFFSET 16'h4070
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_LRCK_ALIGNMENT_BYTE_OFFSET 16'h4080
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_WIDTH 8
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_MASK 8'hff
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_1 8
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_2 16
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_3 24
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_4 32
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_5 40
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_6 48
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_7 56
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_8 64
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_9 72
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_10 80
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_11 88
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_12 96
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_13 104
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_14 112
`define BLOCK_EA_I2S_IN_I2S_INDEX_BIT_OFFSET_15 120
`define BLOCK_EA_I2S_IN_I2S_INDEX_BYTE_WIDTH 16
`define BLOCK_EA_I2S_IN_I2S_INDEX_BYTE_SIZE 16
`define BLOCK_EA_I2S_IN_I2S_INDEX_BYTE_OFFSET 16'h4090
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_WIDTH 32
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_MASK 32'hffffffff
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_1 32
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_2 64
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_3 96
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_4 128
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_5 160
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_6 192
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_7 224
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_8 256
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_9 288
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_10 320
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_11 352
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_12 384
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_13 416
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_14 448
`define BLOCK_EA_I2S_IN_FRAME_NUM_BIT_OFFSET_15 480
`define BLOCK_EA_I2S_IN_FRAME_NUM_BYTE_WIDTH 64
`define BLOCK_EA_I2S_IN_FRAME_NUM_BYTE_SIZE 64
`define BLOCK_EA_I2S_IN_FRAME_NUM_BYTE_OFFSET 16'h4100
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_WIDTH 32
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_MASK 32'hffffffff
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_0 0
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_1 32
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_2 64
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_3 96
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_4 128
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_5 160
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_6 192
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_7 224
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_8 256
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_9 288
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_10 320
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_11 352
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_12 384
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_13 416
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_14 448
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BIT_OFFSET_15 480
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BYTE_WIDTH 64
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BYTE_SIZE 64
`define BLOCK_EA_I2S_IN_BCLK_FREQ_BYTE_OFFSET 16'h4300
`endif
